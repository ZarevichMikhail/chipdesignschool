module top(
    input clk,
    input a,
    input b,
    output q
)


endmodule









