
// Модуль и его название
// top - Название главного модуля в иерархии
module top(

    // входные и выходные сигналы
    input clk,
    input a, // входные и выходные порты могут быть многоразрядными шинами
    input b,
    output q,

    // Для мультиплексора

    input D0,
    input D1,
    input S,
    output Y 

);

// Объявление шины
logic [3:0] c;
logic [8:0] d;

// Присвоить значение можно только в output сигнал
assign q = d[0] // можно присвоить нужный бит
assign q= [4:1] // присваивание диапазона бит
assign q = d[c]; // можно назначить номер бита, определяемый шиной



wire [10:0] a = 7;  // 32-х битное десятичное число, которое будет обрезано
wire [10:0] b = 'd7;  // 11-ти битное десятичное число
wire [10:0] b = 11'd7;  // 11-ти битное десятичное число
wire [3: 0] c = 4'b0101;  // 4-х битное двоичное число
wire [7: 0] d = 8'h7B;  / 8-ми битное шестнадцатеричное число 7B
wire [47:0] e = 48'hEFCA7ED98F;  // 48-ми битное шестнадцатеричное число EFCA7ED98F
wire signed [10:0] b = -11'd7;  // 11-ти битное отрицательное десятичное число



logic [1:0] c; // многобайстный сигнал

assign c = {a,b}; // Конкатенация 


assign Y = S ? D1:D0;




// Конец модуля
endmodule


