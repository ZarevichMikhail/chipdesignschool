`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

    // assign led        = '0;
       //assign abcdefgh   = '0;
       //assign digit      = '0;
       assign red        = '0;
       assign green      = '0;
       assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    logic [31:0] cnt;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            cnt <= '0;
        else
            cnt <= cnt + 1'd1;

    wire enable = (cnt [22:0] == '0);

    //------------------------------------------------------------------------

    wire button_on = | key;

    logic [w_led - 1:0] shift_reg;


    // Задание 1
    /*
    always_ff @ (posedge clk or posedge rst)
        if (rst)
            shift_reg <= '1;
        else if (enable)
            // Светодиоды мигают от 1 до 4
            //shift_reg <= { button_on, shift_reg [w_led - 1:1] };

            // Светодиоды мигают в противоположном направлении. 
            shift_reg <= { shift_reg [w_led - 2:0], button_on };
    assign led = shift_reg;
    */
    // Exercise 1: Make the light move in the opposite direction.




    // Exercise 2: Make the light moving in a loop.
    // Use another key to reset the moving lights back to no lights.

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            //shift_reg <= '1;
            shift_reg <= 'd1;

        else if (key[0])
            shift_reg <='0; // сброс в no lights
        
        // Снова запускает счётчик 
        else if (key[1])
            shift_reg <= 'd1;


        else if (enable)
            // Эта строка реализует циклический сдвиг ВЛЕВО
            // Бит [7] (самый левый) -> в бит [0] (самый правый)
            shift_reg <= { shift_reg[w_led - 2:0], shift_reg[w_led - 1] };


    assign led = shift_reg;
    

    // Exercise 3: Display the state of the shift register
    // on a seven-segment display, moving the light in a circle.

    /*
    always_ff @ (posedge clk or posedge rst)
        if (rst)
            shift_reg <= '1;
        else if (enable)
            // Светодиоды мигают от 1 до 4
            //shift_reg <= { button_on, shift_reg [w_led - 1:1] };

            // Светодиоды мигают в противоположном направлении. 
            shift_reg <= { shift_reg [w_led - 2:0], button_on };
    assign led = shift_reg;

    //------------------------------------------------------------------------
    // ЗАДАНИЕ 3: Счётчик 0-3 на 7-сегментном индикаторе
    //------------------------------------------------------------------------

    // 1. Определим константы для цифр "0", "1", "2", "3" и "Пусто"
    //    Предполагаем, что индикатор с ОБЩИМ АНОДОМ ('0' = сегмент горит)
    localparam PATTERN_0     = 8'b10000001; // Узор для "0"
    localparam PATTERN_1     = 8'b11111001; // Узор для "1"
    localparam PATTERN_2     = 8'b01001001; // Узор для "2"
    localparam PATTERN_3     = 8'b01100001; // Узор для "3"
    localparam PATTERN_BLANK = 8'b11111111; // Все сегменты выключены

    // 2. Создадим новый 2-битный счётчик (00 -> 01 -> 10 -> 11)
    //    Он будет увеличиваться по тому же сигналу 'enable', что и бегущий огонек.
    logic [1:0] count_2bit;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            count_2bit <= '0;
        else if (enable) // Используем тот же медленный 'enable'
            count_2bit <= count_2bit + 1'd1;

    // 3. Логика динамической индикации (мультиплексирование)
    //    Используем быстрый сканер, как в прошлый раз
    logic [2:0] digit_sel;
    assign digit_sel = cnt[15:13]; // 3-битный селектор (000...111)

    // 4. Логика выбора узора
    //    Нам нужно отобразить значение 'count_2bit' (0, 1, 2 или 3)
    //    Мы будем показывать его только на одном, самом правом
    //    индикаторе (digit[0]).
    logic [7:0] current_pattern;

    always_comb
    begin
        // Сначала решим, какой узор (0, 1, 2 или 3) нам нужен
        case (count_2bit)
            2'd0:    current_pattern = PATTERN_0;
            2'd1:    current_pattern = PATTERN_1;
            2'd2:    current_pattern = PATTERN_2;
            2'd3:    current_pattern = PATTERN_3;
            default: current_pattern = PATTERN_BLANK;
        endcase

        // Теперь решим, где (на какой цифре) его показать
        if (digit_sel == 3'd0) // Показываем только на digit[0]
            abcdefgh = current_pattern;
        else
            abcdefgh = PATTERN_BLANK; // Остальные цифры выключены
    end

    // 5. Активируем НУЖНУЮ цифру (дешифратор с активным нулем)
    assign digit = ~(1'b1 << digit_sel);
    */



endmodule
